module motoro3_line_calc_parameter(
    lcStep                   
);

input   wire    [3:0]       lcStep           ;	


endmodule
