module motoro3_line_calc_parameter(
    lSetp                   
);

input   wire    [3:0]       lSetp           ;	


endmodule
