module clk50mhz_to_clk10mhz(
    clk10mhz,
    nRst,
    clk50mhz

);

output  wire                clk10mhz ;	
input   wire                nRst;		
input   wire                clk50mhz;

endmodule
